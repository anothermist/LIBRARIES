// *****************************************************
// AVR address constants (localparams)
//  for registers used by Xcelerator Blocks (XBs) 
// *****************************************************

// Register defines needed for XLR8Float are included as 
// default in the avr_adr_pack.vh located in 
// ../../../XLR8Core/extras/rtl/

